<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 19.0.0, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<!DOCTYPE svg PUBLIC "-//W3C//DTD SVG 1.1//EN" "http://www.w3.org/Graphics/SVG/1.1/DTD/svg11.dtd">
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="0 0 306.1 113.8" style="enable-background:new 0 0 306.1 113.8;" xml:space="preserve">
<style type="text/css">
	.st0{fill:#D0123B;}
	.st1{fill:#D0133C;}
	.st2{fill:#CF113A;}
	.st3{fill:#D0123C;}
	.st4{fill:#CF113B;}
	.st5{fill:#D0153E;}
	.st6{fill:#D0143D;}
</style>
<g>
	<path class="st0" d="M201.8,114c-1.7-1.1-3.4-2.2-4.4-4.2c-1.8,2-3.9,3.2-6.5,3.5c-2.8,0.4-5.7,0.4-8.4-0.7
		c-4.1-1.6-6.3-5.1-6.2-10.1c0.1-6.2,3.6-10,10.3-11.2c2.5-0.4,5-0.6,7.5-0.5c0.7,0,1-0.1,0.9-0.9c-0.1-0.9,0-1.8-0.2-2.6
		c-0.4-2.1-1.4-2.9-3.5-3c-3.5-0.1-6.7,1.1-9.6,2.9c-1.1,0.7-1.5,0.5-2-0.6c-0.7-1.4-1.5-2.7-2.3-4.1c-0.2-0.4-0.3-0.7,0.2-1
		c5.8-3.5,11.9-5.7,18.8-4.2c4.9,1.1,7.4,4,7.5,9c0.1,4.8,0.1,9.6,0,14.4c0,2.8,0.5,5.4,3,7.2c0.6,0.4,0.2,0.7-0.1,1
		c-1.3,1.4-2.6,2.8-3.9,4.2c-0.2,0.2-0.5,0.3-0.4,0.7C202.3,114,202.1,114,201.8,114z M195,101c0-1.1,0-2.2,0-3.4
		c0-0.6-0.2-0.8-0.7-0.8c-1.4,0-2.9,0.1-4.3,0.4c-3.5,0.9-5,4.7-3.2,7.8c0.8,1.3,2,1.9,3.5,1.9c1.2,0,2.3-0.4,3.4-1
		c0.9-0.6,1.5-1.2,1.3-2.4C194.9,102.7,195,101.9,195,101z"/>
	<path class="st1" d="M306.1,48.9c0,0-1.9,0.7-2.7,0.9c-3.3,0.9-6.5,1.2-9.8,0c-3.8-1.4-5.2-3.8-5.3-8.6c0-6.1,0-18.4,0-18.4l0-1.3
		l-3.5,0V15l3.5,0V7.3l9.1-1.5l0,9.5c0,0,5.3,0,7.4,0c0.6,0,0.8,0.2,0.5,0.7c-0.6,1.6-1.3,3.3-1.9,4.9c-0.2,0.6-0.5,0.7-1.1,0.7
		c-1.4,0-2.8,0-4.2,0c-0.5,0-0.8,0.1-0.7,0.6c0.1,6.1-0.1,12.2,0.1,18.4c0.1,3.1,1.8,4.2,5.1,3.5c2-0.4,2-0.4,2-0.4L306.1,48.9z"/>
	<path class="st2" d="M18.8,57.6C12.9,51.7,7,45.9,1.1,40.1c-0.4-0.4-0.6-0.9-0.6-1.5c0-11.5,0-23,0-34.5C0.5,3.2,0.7,3,1.5,3
		c11.6,0,23.2,0,34.8,0c0.7,0,1.1,0.3,1.6,0.7c5.6,5.6,11.3,11.2,16.9,16.8c0.6,0.6,1,0.7,1.7,0C62,14.9,67.7,9.4,73.2,3.8
		c0.6-0.6,1.1-0.9,2-0.9c11.4,0,22.9,0,34.3,0c0.9,0,1.1,0.3,1.1,1.2c0,11.5,0,23,0,34.5c0,0.7-0.2,1.2-0.7,1.7
		c-5.6,5.5-11.1,11-16.6,16.5c-0.3,0.3-0.6,0.6-0.9,1c-0.1,0-0.1,0-0.2,0c-0.3-0.8-1.1-1.2-1.7-1.8C79.3,44.9,68.1,33.8,56.9,22.7
		c-1.3-1.3-1.3-1.3-2.6,0c-8.8,8.8-17.7,17.6-26.5,26.4c-2.9,2.9-5.8,5.7-8.7,8.5C18.9,57.6,18.9,57.6,18.8,57.6z"/>
	<path class="st2" d="M92.2,57.8c0.1,0,0.1,0,0.2,0c0,0,0,0,0,0c0.1,0.1,0.2,0.2,0.3,0.3c3.8,3.7,7.5,7.4,11.3,11.1
		c2,2,4.1,4.1,6.1,6.1c0.4,0.4,0.5,0.7,0.5,1.3c0,11.7,0,23.4,0,35c0,0.8-0.2,1-1,1c-11.6,0-23.1,0-34.7,0c-0.7,0-1.1-0.3-1.5-0.7
		c-5.6-5.6-11.2-11.1-16.7-16.7c-0.8-0.9-1.2-0.7-2,0c-5.5,5.5-11,10.9-16.5,16.4c-0.7,0.7-1.4,0.9-2.3,0.9c-11.4,0-22.7,0-34.1,0
		c-1.1,0-1.3-0.3-1.3-1.3c0-11.4,0-22.7,0-34.1c0-0.8,0.3-1.4,0.8-2c5.6-5.5,11.1-11,16.7-16.6c0.3-0.3,0.7-0.5,0.8-1
		c0.1,0,0.2,0,0.2,0c0.2,0.8,1,1.1,1.5,1.6c8.5,8.5,17,16.9,25.5,25.4c3,2.9,5.9,5.9,8.8,8.8c0.6,0.6,0.9,0.7,1.5,0
		c1.1-1.2,2.3-2.3,3.5-3.5C70.6,79.2,81.4,68.5,92.2,57.8z"/>
	<path class="st3" d="M137.8,25.8c0,7.6,0,15.1,0,22.7c0,1-0.3,1.3-1.3,1.2c-2.5-0.1-5,0-7.4,0c-0.7,0-0.9-0.2-0.9-0.9
		c0-15,0-29.9,0-44.9c0-0.9,0.4-1,1.1-1c2.4,0,4.9,0.1,7.3,0c1,0,1.3,0.2,1.3,1.2c0,6.2,0,12.5,0,18.7c0,0.3,0,0.6,0,0.9
		c0.5-0.2,0.7-0.7,0.9-1.1c3.9-6.2,7.8-12.4,11.7-18.7c0.5-0.8,1-1.1,2-1.1c3.2,0.1,6.5,0,9.7,0c0.1,0.5-0.2,0.7-0.4,1
		c-4.4,6.4-8.7,12.9-13.1,19.3c-0.7,1-0.7,1.6-0.1,2.6c5,7.5,9.8,15.1,14.7,22.7c0.2,0.3,0.5,0.6,0.5,1.1c-3.8,0-7.6,0-11.4,0
		c-0.6,0-0.8-0.5-1-0.9c-4.3-7.3-8.6-14.7-12.9-22C138.4,26.5,138.3,26.1,137.8,25.8z"/>
	<path class="st3" d="M237.4,18.2c-0.2-2.5,1.2-3,3-3.1c1.2-0.1,2.3-0.3,3.4-0.5c0.6-0.1,0.9,0,0.9,0.7c0,5.3-0.1,10.6-0.1,15.9
		c0,6.2,0,12.4,0,18.6c0,1.4-0.1,2.9-0.3,4.3c-0.9,5.5-3.4,8.2-8.9,9.5c-6.5,1.5-12.7,0.4-18.6-2.5c-0.6-0.3-0.6-0.7-0.4-1.2
		c0.6-1.5,1.1-3,1.6-4.5c0.2-0.8,0.4-1,1.3-0.6c3.3,1.6,6.8,2.7,10.5,2.5c0.8,0,1.7-0.1,2.5-0.3c2-0.4,3.2-1.7,3.5-3.7
		c0.1-0.7,0.2-1.5,0.2-2.3c0-1.3,0-2.5,0-4c-1.5,1.6-3.2,2.5-5.1,2.9c-4.7,0.9-11.6-0.6-14.3-8c-2.5-6.8-2.2-13.6,0.9-20.1
		c2.7-5.7,9.2-8.5,14.9-6.7C234.3,15.7,235.8,16.7,237.4,18.2z M236.1,31.4c0-2.4,0-4.4,0-6.4c0-0.4,0-0.9-0.4-1.2
		c-1.8-1.6-3.9-2.1-6.2-1.6c-2.2,0.5-3.2,2.1-3.7,4.2c-0.9,4.2-0.9,8.4,0,12.6c0.6,3,2.5,4.3,5.7,4.1c2.5-0.1,4-1.8,4.4-4.7
		C236.3,35.9,236,33.5,236.1,31.4z"/>
	<path class="st1" d="M260.6,18.3c3.8-3.7,8.1-4.6,13-3.6c4.4,1,6.6,3.9,6.6,9c0.1,8.4,0,16.7,0,25.1c0,0.8-0.3,0.9-1,0.9
		c-2.3,0-4.6-0.1-6.8,0c-0.9,0-1.1-0.3-1.1-1.1c0-7.2,0-14.4,0-21.6c0-0.3,0-0.6,0-1c-0.1-3.3-1.7-4.6-5-3.9c-3.7,0.8-5.5,3-5.6,7.2
		c-0.1,6.3-0.1,12.6,0,18.9c0,1-0.2,1.4-1.3,1.4c-2.4-0.1-4.7-0.1-7.1,0c-0.7,0-1-0.2-1-0.9c0-14.8,0-29.6,0-44.4
		c0-0.6,0.1-0.9,0.7-1c2.6-0.4,5.3-0.8,7.9-1.3c0.8-0.1,0.7,0.4,0.7,0.9c0,4.9,0,9.8-0.1,14.8C260.6,17.9,260.6,18,260.6,18.3z"/>
	<path class="st4" d="M254.9,93.3c0,2.4,0,4.8,0,7.2c0,3.6,0,7.2,0,10.8c0,0.8-0.1,1.1-1,1.1c-2.4-0.1-4.9,0-7.3,0
		c-0.7,0-0.9-0.2-0.9-0.9c0-14.7,0-29.4,0-44.1c0-0.6,0.2-0.9,0.8-1c2.6-0.4,5.1-0.8,7.7-1.2c0.9-0.1,0.7,0.4,0.7,0.9
		c0,4.3,0,8.6,0,13c0,4.4,0,8.8,0,13.3c0.5-0.2,0.6-0.6,0.8-0.9c2.5-4.2,5.1-8.4,7.6-12.6c0.4-0.6,0.8-0.9,1.5-0.9
		c3.3,0,6.6,0,10.1,0c-0.8,1-1.4,1.8-2,2.6c-2.8,3.7-5.7,7.3-8.5,11c-0.6,0.7-0.5,1.1,0,1.8c4.3,6.3,8.6,12.6,12.9,18.9
		c-0.2,0.4-0.6,0.2-0.9,0.2c-2.9,0-5.8,0-8.6,0c-0.8,0-1.3-0.2-1.7-0.9c-3.5-5.8-7-11.5-10.5-17.3C255.5,93.8,255.4,93.4,254.9,93.3
		z"/>
	<path class="st5" d="M219.8,81.8c3-3.2,6.4-4.7,10.6-4.5c5.3,0.2,8.5,3.3,8.5,8.6c0.1,8.5,0,17,0,25.6c0,0.8-0.2,0.9-1,0.9
		c-2.3,0-4.6-0.1-7,0c-0.9,0-1-0.3-1-1.1c0-7,0-14.1,0-21.1c0-0.6,0-1.3-0.1-1.9c-0.3-2.8-1.9-3.9-4.6-3.1c-2.6,0.8-4.4,2.9-4.5,5.7
		c-0.1,3.6-0.1,7.1-0.1,10.7c0,3.2,0,6.5,0,9.7c0,0.8-0.1,1.1-1,1.1c-2.4-0.1-4.8,0-7.2,0c-0.7,0-1-0.2-1-0.9c0-10.6,0-21.3,0-31.9
		c0-0.7,0.1-1,0.9-1.1c2.1-0.3,4.1-0.6,6.1-1c0.6-0.1,0.8,0.1,0.8,0.7C219.5,79.2,219.6,80.4,219.8,81.8z"/>
	<path class="st1" d="M175,19.2c0.3-0.4,0.5-0.8,0.8-1.1c3.3-3,7.3-4.1,11.7-3.1c4.2,1,6.3,3.7,6.3,8.3c0.1,8.5,0,17,0,25.6
		c0,0.7-0.2,0.9-1,0.9c-2.3,0-4.6-0.1-6.8,0c-0.9,0-1.1-0.2-1.1-1.1c0-6.9,0-13.8,0-20.8c0-0.9-0.1-1.8-0.2-2.6
		c-0.3-2.4-1.7-3.4-4.1-2.8c-2.9,0.6-4.9,3-5,6.1c-0.1,4.6-0.1,9.3-0.1,13.9c0,2.1,0,4.2,0,6.4c0,0.7-0.2,1-0.9,0.9
		c-2.4,0-4.9-0.1-7.3,0c-0.8,0-1-0.3-1-1c0-4,0-8,0-12c0-6.4,0-12.9,0-19.3c0-1.1,0.2-1.6,1.4-1.7c1.9-0.2,3.7-0.6,5.6-0.9
		c0.6-0.1,0.9,0,1,0.7c0.1,1.1,0.3,2.3,0.5,3.4C174.8,19.1,174.9,19.1,175,19.2z"/>
	<path class="st1" d="M128.1,88.9c0-7.4,0-14.8,0-22.2c0-0.9,0.2-1.2,1.2-1.2c7.7,0,15.4,0,23.2,0c0.9,0,1.2,0.1,1,1.2
		c-0.4,1.8-0.6,3.5-0.8,5.3c-0.1,0.9-0.5,1.1-1.3,1.1c-4.3,0-8.6,0-12.8,0c-0.8,0-1.1,0.2-1.1,1.1c0,2.9,0,5.8,0,8.8
		c0,0.8,0.2,1.1,1.1,1.1c3.3,0,6.6,0,10,0c0.8,0,1.1,0.2,1.1,1.1c-0.1,1.9-0.1,3.8,0,5.6c0,0.8-0.2,1-1,1c-3.3,0-6.6,0-9.8,0
		c-1,0-1.3,0.2-1.3,1.2c0.1,6.1,0,12.2,0,18.4c0,0.9-0.2,1.2-1.1,1.1c-2.4-0.1-4.7-0.1-7.1,0c-1,0-1.1-0.4-1.1-1.2
		C128.1,103.7,128.1,96.3,128.1,88.9z"/>
	<path class="st6" d="M163.1,82.2c1.1-1.4,2.2-2.6,3.5-3.5c2.2-1.6,4.6-2.1,7.3-1.3c0.6,0.2,0.9,0.4,0.6,1.2
		c-0.7,2.1-1.2,4.2-1.8,6.3c-0.2,0.7-0.4,0.9-1.1,0.6c-0.9-0.4-1.8-0.5-2.8-0.4c-2.9,0.3-4.5,1.9-4.7,4.8c-0.2,3.2-0.1,6.5-0.1,9.7
		c0,3.9,0,7.8,0,11.6c0,0.9-0.2,1.1-1.1,1.1c-2.4-0.1-4.7,0-7.1,0c-0.7,0-1-0.1-1-1c0-10.5,0-21,0-31.6c0-0.7,0.2-1,1-1.1
		c1.8-0.2,3.6-0.6,5.4-0.9c0.8-0.1,1.2,0,1.3,0.9C162.6,79.8,162.9,80.8,163.1,82.2z"/>
	<path class="st5" d="M209.9,32.1c0,5.5,0,10.9,0,16.4c0,1-0.3,1.2-1.2,1.2c-2.3-0.1-4.6-0.1-7,0c-0.8,0-1.1-0.1-1.1-1
		c0-10.6,0-21.2,0-31.8c0-0.7,0.1-1,0.9-1.1c2.4-0.3,4.8-0.7,7.2-1.2c0.8-0.1,1.1,0.1,1.1,0.9C209.9,21.1,209.9,26.6,209.9,32.1z"/>
	<path class="st2" d="M92.7,58.1c-0.1-0.1-0.2-0.2-0.3-0.3C92.5,57.9,92.6,58,92.7,58.1z"/>
</g>
<circle class="st1" cx="205.3" cy="5.9" r="5.7"/>
</svg>
